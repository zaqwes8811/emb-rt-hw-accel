
module ni2 (
	clk_clk,
	pio_external_connection_export);	

	input		clk_clk;
	output	[7:0]	pio_external_connection_export;
endmodule
