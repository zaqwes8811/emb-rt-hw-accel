`timescale 10ns/1ps


// fixme: memory access unregular - сделать пока просто, с поворотом
//  потом думать об оптимизации - пока сложно представить

// rect:
// https://www.researchgate.net/profile/Ratiba_Fellag/publication/273348053_Survey_on_Image_Rectification_on_FPGA/links/54ff043f0cf2672e2240f3a5.pdf

module homography_warp_tb;

endmodule