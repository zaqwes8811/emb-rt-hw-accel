`timescale 10ns/1ps


// fixme: memory access unregular - сделать пока просто, с поворотом
//  потом думать об оптимизации - пока сложно представить

module homography_warp_tb;

endmodule